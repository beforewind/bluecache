import ClientServer::*;
interface Server#(


interface LockServer#(numeric type numServers);
   interface Vector#(numServers, 
